module KeyboardCtrl#(
   parameter SYSCLK_FREQUENCY_HZ = 100000000
)(
    output reg [7:0] key_in,
    output reg is_extend,
    output reg is_break,
		output reg valid,
    output err,
    inout PS2_DATA,
    inout PS2_CLK,
    input rst,
    input clk
);
//////////////////////////////////////////////////////////
// This Keyboard  Controller do not support lock LED control
//////////////////////////////////////////////////////////

  parameter RESET          = 3'd0;
	parameter SEND_CMD       = 3'd1;
	parameter WAIT_ACK       = 3'd2;
  parameter WAIT_KEYIN     = 3'd3;
	parameter GET_BREAK      = 3'd4;
	parameter GET_EXTEND     = 3'd5;
	parameter RESET_WAIT_BAT = 3'd6;
    
  parameter CMD_RESET           = 8'hFF; 
  parameter CMD_SET_STATUS_LEDS = 8'hED;
	parameter RSP_ACK             = 8'hFA;
	parameter RSP_BAT_PASS        = 8'hAA;
    
  parameter BREAK_CODE  = 8'hF0;
  parameter EXTEND_CODE = 8'hE0;
  parameter CAPS_LOCK   = 8'h58;
  parameter NUM_LOCK    = 8'h77;
  parameter SCR_LOCK    = 8'h7E;
    
  wire [7:0] rx_data;
	wire rx_valid;
	wire busy;
	
	reg [7:0] tx_data;
	reg tx_valid;
	reg [2:0] state;
	reg [2:0] lock_status;
	
	always @ (posedge clk, posedge rst)
	  if(rst)
	    key_in <= 0;
	  else if(rx_valid)
	    key_in <= rx_data;
	  else
	    key_in <= key_in;
	
	always @ (posedge clk, posedge rst) begin
	  if (rst) begin
	    state <= RESET;
      is_extend <= 1'b0;
      is_break <= 1'b1;
			valid <= 1'b0;
			lock_status <= 3'b0;
			tx_data <= 8'h00;
			tx_valid <= 1'b0;
	  end else begin
	    is_extend <= 1'b0;
	    is_break <= 1'b0;
	    valid <= 1'b0;
	    lock_status <= lock_status;
	    tx_data <= tx_data;
	    tx_valid <= 1'b0;
	    case (state)
			RESET: begin
				is_extend <= 1'b0;
				is_break <= 1'b1;
				valid <= 1'b0;
				lock_status <= 3'b0;
				tx_data <= CMD_RESET;
				tx_valid <= 1'b0;
				state <= SEND_CMD;
				end
		  
		  SEND_CMD: begin
		    if (busy == 1'b0) begin
			    tx_valid <= 1'b1;
					state <= WAIT_ACK;
			  end else begin
			    tx_valid <= 1'b0;
					state <= SEND_CMD;
		    end
		  end
	      
		  WAIT_ACK: begin
				if(rx_valid == 1'b1) begin
					if (rx_data == RSP_ACK && tx_data == CMD_RESET) begin
					state <= RESET_WAIT_BAT;
					end else if (rx_data == RSP_ACK && tx_data == CMD_SET_STATUS_LEDS) begin
						tx_data <= {5'b00000, lock_status};
						state <= SEND_CMD;
					end else begin
						state <= WAIT_KEYIN;
					end
				end else if (err == 1'b1) begin
					state <= RESET;
				end else begin
					state <= WAIT_ACK;
				end
		  end
			
		  WAIT_KEYIN: begin
				if (rx_valid == 1'b1 && rx_data == BREAK_CODE) begin
					state <= GET_BREAK;
				end else if (rx_valid == 1'b1 && rx_data == EXTEND_CODE) begin
					state <= GET_EXTEND;
				end else if (rx_valid == 1'b1) begin
					state <= WAIT_KEYIN;
					valid <= 1'b1;
				end else if (err == 1'b1) begin
					state <= RESET;
				end else begin
					state <= WAIT_KEYIN;
				end
			end
		    
		  GET_BREAK: begin
		    is_extend <= is_extend;
		    if (rx_valid == 1'b1) begin
					state <= WAIT_KEYIN;
					valid <= 1'b1;
					is_break <= 1'b1;
			  end else if (err == 1'b1) begin
			    state <= RESET;
			  end else begin
			    state <= GET_BREAK;
			  end
		  end
			
		  GET_EXTEND: begin
		    if (rx_valid == 1'b1 && rx_data == BREAK_CODE) begin
		      state <= GET_BREAK;
		      is_extend <= 1'b1;
		    end else if (rx_valid == 1'b1) begin
		      state <= WAIT_KEYIN;
          valid <= 1'b1;
		      is_extend <= 1'b1;
			  end else if (err == 1'b1) begin
			  	state <= RESET;
		    end else begin
		      state <= GET_EXTEND;
		    end
		  end
			
		  RESET_WAIT_BAT: begin
		    if (rx_valid == 1'b1 && rx_data == RSP_BAT_PASS) begin
			    state <= WAIT_KEYIN;
			  end else if (rx_valid == 1'b1) begin
			    state <= RESET;
			  end else if (err == 1'b1) begin
			    state <= RESET;
			  end else begin
			    state <= RESET_WAIT_BAT;
			  end
		  end

		  default: begin
		    state <= RESET;
		    valid <= 1'b0;
		  end
		endcase
	  end
	end
	
    Ps2Interface #(
      .SYSCLK_FREQUENCY_HZ(SYSCLK_FREQUENCY_HZ)
    ) Ps2Interface_i(
      .ps2_clk(PS2_CLK),
      .ps2_data(PS2_DATA),
      
      .clk(clk),
      .rst(rst),
      
      .tx_data(tx_data),
      .tx_valid(tx_valid),
      
      .rx_data(rx_data),
      .rx_valid(rx_valid),
      
      .busy(busy),
      .err(err)
    );
        
endmodule
